typedef uvm_sequencer #(apb_tx)apb_sqr;
