`include "uvm_pkg.sv"
import uvm_pkg::*;

`include "mem.v"
`include "apb_common.sv"
`include "apb_intrf.sv"
`include "apb_tx.sv"
`include "apb_seq_lib.sv"
`include "apb_sqr.sv"
`include "apb_drv.sv"
`include "apb_mon.sv"
`include "apb_cov.sv"
`include "apb_agent.sv"
`include "apb_sbd.sv"
`include "apb_env.sv"
`include "apb_base_test.sv"
`include "top.sv"
